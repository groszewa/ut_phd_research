parameter DATA_WIDTH  = {{ data.get('data_width')    }};
parameter NUM_INPUTS  = {{ data.get('num_inputs')    }};
parameter WXIP1       = {{ data.get('wxip1')         }};
parameter MIN_CYC_DSC = {{ data.get('min_cycle_dsc') }};

