parameter DATA_WIDTH = 6;
parameter NUM_INPUTS = 2;
