parameter DATA_WIDTH = 8;
parameter NUM_INPUTS = 2;
parameter WXIP1 = 17;
parameter MIN_CYC_DSC = 256;

