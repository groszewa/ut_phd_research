parameter DATA_WIDTH = 6;
parameter NUM_INPUTS = 2;
parameter WXIP1 = 13;
parameter MIN_CYC_DSC = 1234;

