`timescale 1 ns / 100 ps


module ms_es_ordered_bs_by4_mul #(parameter DATA_WIDTH=5, parameter NUM_INPUTS=2, parameter WXIP1=1) (
	clk,
	rst,
	en,
	bin_data_in,
	bin_data_out,
	done);

	input  [DATA_WIDTH-1:0] bin_data_in [NUM_INPUTS-1:0];
	input                   clk,rst,en;

	output [WXIP1-1:0] bin_data_out;
	output                               done;
	
	wire [NUM_INPUTS-1:0] sng_ov;
    wire [3:0]             bs_data_in [NUM_INPUTS-1:0];
   
   
	wire [4**(NUM_INPUTS)-1:0] bs_data_out;
	wire dummy_ov;
   
	genvar i;
	generate
		for(i=0;i<NUM_INPUTS;i++) begin
			if(i==0) begin
				sng_dsc_ms_max #(.WIDTH(DATA_WIDTH), .NUM_INPUTS(NUM_INPUTS), .STRIDE(4)) sng (
					.clk(clk),
					.rst(rst),
					.en(en),
					.bin_in(bin_data_in),
					.sn_out(bs_data_in[0]),
					.ctr_overflow(sng_ov[0]));
            end
			if (i==NUM_INPUTS-1) begin
				sng_dsc_ms_min #(.WIDTH(DATA_WIDTH), .NUM_INPUTS(NUM_INPUTS), .STRIDE(4)) sng (
					.clk(sng_ov[i-1]),
					.rst(rst),
					.en(en),
					.bin_in(bin_data_in),
					.sn_out(bs_data_in[i]),
					.ctr_overflow(sng_ov[i]));
			end
            if (NUM_INPUTS==3) begin
               if (i==1) begin
 				sng_dsc_ms_mid_of3 #(.WIDTH(DATA_WIDTH), .NUM_INPUTS(NUM_INPUTS), .STRIDE(4)) sng (
					.clk(sng_ov[i-1]),
					.rst(rst),
					.en(en),
					.bin_in(bin_data_in),
					.sn_out(bs_data_in[i]),
					.ctr_overflow(sng_ov[i]));                 
               end
            end
            if (NUM_INPUTS==4) begin
               if (i==1) begin
  				  sng_dsc_ms_second_largest_of4 #(.WIDTH(DATA_WIDTH), .NUM_INPUTS(NUM_INPUTS), .STRIDE(4)) sng (
					  .clk(sng_ov[i-1]),
					  .rst(rst),
					  .en(en),
					  .bin_in(bin_data_in),
					  .sn_out(bs_data_in[i]),
					  .ctr_overflow(sng_ov[i]));                 
               end
               if (i==2) begin
  				  sng_dsc_ms_second_smallest_of4 #(.WIDTH(DATA_WIDTH), .NUM_INPUTS(NUM_INPUTS), .STRIDE(4)) sng (
					  .clk(sng_ov[i-1]),
					  .rst(rst),
					  .en(en),
					  .bin_in(bin_data_in),
					  .sn_out(bs_data_in[i]),
					  .ctr_overflow(sng_ov[i]));                                   
               end
            end
            if (NUM_INPUTS==5) begin
               if (i==1) begin
   				  sng_dsc_ms_second_largest_of5 #(.WIDTH(DATA_WIDTH), .NUM_INPUTS(NUM_INPUTS), .STRIDE(4)) sng (
					  .clk(sng_ov[i-1]),
					  .rst(rst),
					  .en(en),
					  .bin_in(bin_data_in),
					  .sn_out(bs_data_in[i]),
					  .ctr_overflow(sng_ov[i]));                                  
               end
               if (i==2) begin
  				  sng_dsc_ms_mid_of5 #(.WIDTH(DATA_WIDTH), .NUM_INPUTS(NUM_INPUTS), .STRIDE(4)) sng (
					  .clk(sng_ov[i-1]),
					  .rst(rst),
					  .en(en),
					  .bin_in(bin_data_in),
					  .sn_out(bs_data_in[i]),
					  .ctr_overflow(sng_ov[i]));                                   
               end
               if (i==3) begin
  				  sng_dsc_ms_second_smallest_of5 #(.WIDTH(DATA_WIDTH), .NUM_INPUTS(NUM_INPUTS), .STRIDE(4)) sng (
					  .clk(sng_ov[i-1]),
					  .rst(rst),
					  .en(en),
					  .bin_in(bin_data_in),
					  .sn_out(bs_data_in[i]),
					  .ctr_overflow(sng_ov[i]));                                   
               end
            end
		end
	endgenerate	


    //FIXME
	//assign bs_data_out = &bs_data_in;
    //multiplier circuit calculates (a0+a1)*(b0+b1)=a0b0+a0b1+a1b0+a1b1
    //genvar j;
    //for(i=0;i<2;i++) begin
    //   for(j=0;j<2;j++) begin
    //      assign bs_data_out[{i,j}] = bs_data_in[0][i] & bs_data_in[1][j];
    //   end
    //end
   if (NUM_INPUTS==2) begin
      assign bs_data_out[0]  = bs_data_in[0][0] & bs_data_in[1][0];
      assign bs_data_out[1]  = bs_data_in[0][0] & bs_data_in[1][1];
      assign bs_data_out[2]  = bs_data_in[0][0] & bs_data_in[1][2];
      assign bs_data_out[3]  = bs_data_in[0][0] & bs_data_in[1][3];
      assign bs_data_out[4]  = bs_data_in[0][1] & bs_data_in[1][0];
      assign bs_data_out[5]  = bs_data_in[0][1] & bs_data_in[1][1];
      assign bs_data_out[6]  = bs_data_in[0][1] & bs_data_in[1][2];
      assign bs_data_out[7]  = bs_data_in[0][1] & bs_data_in[1][3];
      assign bs_data_out[8]  = bs_data_in[0][2] & bs_data_in[1][0];
      assign bs_data_out[9]  = bs_data_in[0][2] & bs_data_in[1][1];
      assign bs_data_out[10] = bs_data_in[0][2] & bs_data_in[1][2];
      assign bs_data_out[11] = bs_data_in[0][2] & bs_data_in[1][3];
      assign bs_data_out[12] = bs_data_in[0][3] & bs_data_in[1][0];
      assign bs_data_out[13] = bs_data_in[0][3] & bs_data_in[1][1];
      assign bs_data_out[14] = bs_data_in[0][3] & bs_data_in[1][2];
      assign bs_data_out[15] = bs_data_in[0][3] & bs_data_in[1][3];
      

      par_acc_16lanes  #(.WIDTH(DATA_WIDTH*NUM_INPUTS)) stoch2bin (
        .clk(clk),
        .rst(rst),                                               
        .data_in(bs_data_out),
        .countval(bin_data_out),
        .overflow(dummy_ov));

   end // if (NUM_INPUTS==2)
   else if (NUM_INPUTS==3) begin //FIXME
      assign bs_data_out[0]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0];
      assign bs_data_out[1]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1];
      assign bs_data_out[2]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2];
      assign bs_data_out[3]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3];
      assign bs_data_out[4]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0];
      assign bs_data_out[5]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1];
      assign bs_data_out[6]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2];
      assign bs_data_out[7]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3];
      assign bs_data_out[8]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0];
      assign bs_data_out[9]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1];
      assign bs_data_out[10] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2];
      assign bs_data_out[11] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3];
      assign bs_data_out[12] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0];
      assign bs_data_out[13] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1];
      assign bs_data_out[14] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2];
      assign bs_data_out[15] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3];
      assign bs_data_out[16] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0];
      assign bs_data_out[17] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1];
      assign bs_data_out[18] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2];
      assign bs_data_out[19] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3];
      assign bs_data_out[20] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0];
      assign bs_data_out[21] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1];
      assign bs_data_out[22] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2];
      assign bs_data_out[23] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3];
      assign bs_data_out[24] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0];
      assign bs_data_out[25] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1];
      assign bs_data_out[26] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2];
      assign bs_data_out[27] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3];
      assign bs_data_out[28] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0];
      assign bs_data_out[29] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1];
      assign bs_data_out[30] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2];
      assign bs_data_out[31] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3];
      assign bs_data_out[32] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0];
      assign bs_data_out[33] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1];
      assign bs_data_out[34] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2];
      assign bs_data_out[35] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3];
      assign bs_data_out[36] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0];
      assign bs_data_out[37] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1];
      assign bs_data_out[38] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2];
      assign bs_data_out[39] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3];
      assign bs_data_out[40] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0];
      assign bs_data_out[41] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1];
      assign bs_data_out[42] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2];
      assign bs_data_out[43] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3];
      assign bs_data_out[44] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0];
      assign bs_data_out[45] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1];
      assign bs_data_out[46] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2];
      assign bs_data_out[47] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3];
      assign bs_data_out[48] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0];
      assign bs_data_out[49] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1];
      assign bs_data_out[50] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2];
      assign bs_data_out[51] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3];
      assign bs_data_out[52] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0];
      assign bs_data_out[53] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1];
      assign bs_data_out[54] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2];
      assign bs_data_out[55] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3];
      assign bs_data_out[56] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0];
      assign bs_data_out[57] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1];
      assign bs_data_out[58] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2];
      assign bs_data_out[59] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3];
      assign bs_data_out[60] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0];
      assign bs_data_out[61] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1];
      assign bs_data_out[62] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2];
      assign bs_data_out[63] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3];
  
      par_acc_64lanes  #(.WIDTH(DATA_WIDTH*NUM_INPUTS)) stoch2bin (
        .clk(clk),
        .rst(rst),                                               
        .data_in(bs_data_out),
        .countval(bin_data_out),
        .overflow(dummy_ov));

   end // if (NUM_INPUTS==3)
   else if (NUM_INPUTS==4) begin //FIXME
      assign bs_data_out[0]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[1]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[2]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[3]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[4]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[5]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[6]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[7]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[8]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[9]   = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[10]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[11]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[12]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[13]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[14]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[15]  = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[16]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[17]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[18]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[19]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[20]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[21]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[22]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[23]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[24]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[25]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[26]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[27]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[28]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[29]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[30]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[31]  = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[32]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[33]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[34]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[35]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[36]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[37]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[38]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[39]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[40]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[41]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[42]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[43]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[44]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[45]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[46]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[47]  = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[48]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[49]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[50]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[51]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[52]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[53]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[54]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[55]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[56]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[57]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[58]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[59]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[60]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[61]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[62]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[63]  = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[64]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[65]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[66]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[67]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[68]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[69]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[70]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[71]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[72]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[73]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[74]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[75]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[76]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[77]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[78]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[79]  = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[80]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[81]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[82]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[83]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[84]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[85]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[86]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[87]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[88]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[89]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[90]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[91]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[92]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[93]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[94]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[95]  = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[96]  = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[97]  = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[98]  = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[99]  = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[100] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[101] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[102] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[103] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[104] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[105] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[106] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[107] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[108] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[109] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[110] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[111] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[112] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[113] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[114] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[115] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[116] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[117] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[118] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[119] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[120] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[121] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[122] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[123] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[124] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[125] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[126] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[127] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[128] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[129] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[130] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[131] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[132] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[133] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[134] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[135] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[136] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[137] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[138] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[139] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[140] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[141] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[142] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[143] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[144] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[145] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[146] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[147] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[148] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[149] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[150] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[151] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[152] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[153] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[154] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[155] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[156] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[157] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[158] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[159] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[160] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[161] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[162] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[163] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[164] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[165] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[166] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[167] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[168] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[169] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[170] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[171] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[172] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[173] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[174] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[175] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[176] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[177] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[178] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[179] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[180] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[181] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[182] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[183] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[184] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[185] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[186] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[187] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[188] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[189] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[190] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[191] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[192] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[193] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[194] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[195] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[196] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[197] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[198] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[199] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[200] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[201] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[202] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[203] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[204] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[205] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[206] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[207] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[208] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[209] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[210] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[211] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[212] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[213] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[214] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[215] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[216] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[217] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[218] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[219] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[220] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[221] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[222] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[223] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[224] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[225] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[226] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[227] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[228] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[229] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[230] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[231] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[232] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[233] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[234] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[235] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[236] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[237] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[238] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[239] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3];
      assign bs_data_out[240] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0];
      assign bs_data_out[241] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1];
      assign bs_data_out[242] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2];
      assign bs_data_out[243] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3];
      assign bs_data_out[244] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0];
      assign bs_data_out[245] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1];
      assign bs_data_out[246] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2];
      assign bs_data_out[247] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3];
      assign bs_data_out[248] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0];
      assign bs_data_out[249] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1];
      assign bs_data_out[250] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2];
      assign bs_data_out[251] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3];
      assign bs_data_out[252] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0];
      assign bs_data_out[253] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1];
      assign bs_data_out[254] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2];
      assign bs_data_out[255] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3];
  
      par_acc_256lanes  #(.WIDTH(DATA_WIDTH*NUM_INPUTS)) stoch2bin (
        .clk(clk),
        .rst(rst),                                               
        .data_in(bs_data_out),
        .countval(bin_data_out),
        .overflow(dummy_ov));

   end // if (NUM_INPUTS==4)
   else if (NUM_INPUTS==5) begin //FIXME
      assign bs_data_out[0] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[1] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[2] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[3] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[4] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[5] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[6] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[7] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[8] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[9] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[10] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[11] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[12] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[13] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[14] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[15] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[16] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[17] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[18] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[19] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[20] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[21] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[22] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[23] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[24] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[25] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[26] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[27] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[28] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[29] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[30] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[31] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[32] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[33] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[34] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[35] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[36] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[37] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[38] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[39] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[40] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[41] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[42] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[43] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[44] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[45] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[46] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[47] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[48] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[49] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[50] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[51] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[52] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[53] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[54] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[55] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[56] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[57] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[58] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[59] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[60] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[61] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[62] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[63] = bs_data_in[0][0] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[64] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[65] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[66] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[67] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[68] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[69] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[70] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[71] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[72] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[73] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[74] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[75] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[76] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[77] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[78] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[79] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[80] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[81] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[82] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[83] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[84] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[85] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[86] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[87] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[88] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[89] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[90] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[91] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[92] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[93] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[94] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[95] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[96] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[97] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[98] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[99] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[100] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[101] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[102] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[103] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[104] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[105] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[106] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[107] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[108] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[109] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[110] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[111] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[112] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[113] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[114] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[115] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[116] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[117] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[118] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[119] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[120] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[121] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[122] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[123] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[124] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[125] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[126] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[127] = bs_data_in[0][0] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[128] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[129] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[130] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[131] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[132] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[133] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[134] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[135] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[136] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[137] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[138] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[139] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[140] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[141] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[142] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[143] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[144] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[145] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[146] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[147] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[148] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[149] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[150] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[151] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[152] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[153] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[154] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[155] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[156] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[157] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[158] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[159] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[160] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[161] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[162] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[163] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[164] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[165] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[166] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[167] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[168] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[169] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[170] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[171] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[172] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[173] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[174] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[175] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[176] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[177] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[178] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[179] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[180] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[181] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[182] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[183] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[184] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[185] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[186] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[187] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[188] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[189] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[190] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[191] = bs_data_in[0][0] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[192] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[193] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[194] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[195] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[196] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[197] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[198] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[199] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[200] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[201] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[202] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[203] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[204] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[205] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[206] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[207] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[208] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[209] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[210] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[211] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[212] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[213] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[214] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[215] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[216] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[217] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[218] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[219] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[220] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[221] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[222] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[223] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[224] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[225] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[226] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[227] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[228] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[229] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[230] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[231] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[232] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[233] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[234] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[235] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[236] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[237] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[238] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[239] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[240] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[241] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[242] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[243] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[244] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[245] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[246] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[247] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[248] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[249] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[250] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[251] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[252] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[253] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[254] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[255] = bs_data_in[0][0] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[256] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[257] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[258] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[259] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[260] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[261] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[262] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[263] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[264] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[265] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[266] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[267] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[268] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[269] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[270] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[271] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[272] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[273] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[274] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[275] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[276] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[277] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[278] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[279] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[280] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[281] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[282] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[283] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[284] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[285] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[286] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[287] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[288] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[289] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[290] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[291] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[292] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[293] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[294] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[295] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[296] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[297] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[298] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[299] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[300] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[301] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[302] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[303] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[304] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[305] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[306] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[307] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[308] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[309] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[310] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[311] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[312] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[313] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[314] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[315] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[316] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[317] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[318] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[319] = bs_data_in[0][1] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[320] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[321] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[322] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[323] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[324] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[325] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[326] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[327] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[328] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[329] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[330] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[331] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[332] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[333] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[334] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[335] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[336] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[337] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[338] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[339] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[340] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[341] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[342] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[343] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[344] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[345] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[346] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[347] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[348] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[349] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[350] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[351] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[352] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[353] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[354] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[355] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[356] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[357] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[358] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[359] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[360] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[361] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[362] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[363] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[364] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[365] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[366] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[367] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[368] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[369] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[370] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[371] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[372] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[373] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[374] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[375] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[376] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[377] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[378] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[379] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[380] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[381] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[382] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[383] = bs_data_in[0][1] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[384] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[385] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[386] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[387] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[388] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[389] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[390] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[391] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[392] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[393] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[394] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[395] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[396] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[397] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[398] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[399] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[400] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[401] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[402] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[403] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[404] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[405] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[406] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[407] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[408] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[409] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[410] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[411] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[412] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[413] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[414] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[415] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[416] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[417] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[418] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[419] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[420] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[421] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[422] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[423] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[424] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[425] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[426] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[427] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[428] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[429] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[430] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[431] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[432] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[433] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[434] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[435] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[436] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[437] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[438] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[439] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[440] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[441] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[442] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[443] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[444] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[445] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[446] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[447] = bs_data_in[0][1] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[448] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[449] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[450] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[451] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[452] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[453] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[454] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[455] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[456] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[457] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[458] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[459] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[460] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[461] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[462] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[463] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[464] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[465] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[466] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[467] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[468] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[469] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[470] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[471] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[472] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[473] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[474] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[475] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[476] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[477] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[478] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[479] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[480] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[481] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[482] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[483] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[484] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[485] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[486] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[487] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[488] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[489] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[490] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[491] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[492] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[493] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[494] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[495] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[496] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[497] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[498] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[499] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[500] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[501] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[502] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[503] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[504] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[505] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[506] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[507] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[508] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[509] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[510] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[511] = bs_data_in[0][1] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[512] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[513] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[514] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[515] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[516] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[517] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[518] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[519] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[520] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[521] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[522] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[523] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[524] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[525] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[526] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[527] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[528] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[529] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[530] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[531] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[532] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[533] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[534] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[535] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[536] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[537] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[538] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[539] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[540] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[541] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[542] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[543] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[544] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[545] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[546] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[547] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[548] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[549] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[550] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[551] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[552] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[553] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[554] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[555] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[556] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[557] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[558] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[559] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[560] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[561] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[562] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[563] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[564] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[565] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[566] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[567] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[568] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[569] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[570] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[571] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[572] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[573] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[574] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[575] = bs_data_in[0][2] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[576] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[577] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[578] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[579] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[580] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[581] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[582] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[583] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[584] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[585] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[586] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[587] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[588] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[589] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[590] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[591] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[592] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[593] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[594] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[595] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[596] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[597] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[598] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[599] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[600] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[601] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[602] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[603] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[604] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[605] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[606] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[607] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[608] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[609] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[610] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[611] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[612] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[613] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[614] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[615] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[616] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[617] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[618] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[619] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[620] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[621] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[622] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[623] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[624] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[625] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[626] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[627] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[628] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[629] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[630] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[631] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[632] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[633] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[634] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[635] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[636] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[637] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[638] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[639] = bs_data_in[0][2] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[640] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[641] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[642] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[643] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[644] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[645] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[646] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[647] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[648] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[649] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[650] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[651] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[652] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[653] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[654] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[655] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[656] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[657] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[658] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[659] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[660] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[661] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[662] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[663] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[664] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[665] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[666] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[667] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[668] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[669] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[670] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[671] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[672] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[673] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[674] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[675] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[676] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[677] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[678] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[679] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[680] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[681] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[682] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[683] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[684] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[685] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[686] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[687] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[688] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[689] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[690] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[691] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[692] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[693] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[694] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[695] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[696] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[697] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[698] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[699] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[700] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[701] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[702] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[703] = bs_data_in[0][2] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[704] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[705] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[706] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[707] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[708] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[709] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[710] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[711] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[712] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[713] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[714] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[715] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[716] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[717] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[718] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[719] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[720] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[721] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[722] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[723] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[724] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[725] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[726] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[727] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[728] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[729] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[730] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[731] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[732] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[733] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[734] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[735] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[736] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[737] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[738] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[739] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[740] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[741] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[742] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[743] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[744] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[745] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[746] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[747] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[748] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[749] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[750] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[751] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[752] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[753] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[754] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[755] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[756] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[757] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[758] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[759] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[760] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[761] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[762] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[763] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[764] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[765] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[766] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[767] = bs_data_in[0][2] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[768] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[769] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[770] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[771] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[772] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[773] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[774] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[775] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[776] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[777] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[778] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[779] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[780] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[781] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[782] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[783] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[784] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[785] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[786] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[787] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[788] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[789] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[790] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[791] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[792] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[793] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[794] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[795] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[796] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[797] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[798] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[799] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[800] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[801] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[802] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[803] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[804] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[805] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[806] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[807] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[808] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[809] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[810] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[811] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[812] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[813] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[814] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[815] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[816] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[817] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[818] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[819] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[820] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[821] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[822] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[823] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[824] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[825] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[826] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[827] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[828] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[829] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[830] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[831] = bs_data_in[0][3] & bs_data_in[1][0] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[832] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[833] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[834] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[835] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[836] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[837] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[838] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[839] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[840] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[841] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[842] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[843] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[844] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[845] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[846] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[847] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[848] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[849] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[850] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[851] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[852] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[853] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[854] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[855] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[856] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[857] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[858] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[859] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[860] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[861] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[862] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[863] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[864] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[865] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[866] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[867] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[868] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[869] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[870] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[871] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[872] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[873] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[874] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[875] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[876] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[877] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[878] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[879] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[880] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[881] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[882] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[883] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[884] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[885] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[886] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[887] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[888] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[889] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[890] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[891] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[892] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[893] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[894] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[895] = bs_data_in[0][3] & bs_data_in[1][1] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[896] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[897] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[898] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[899] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[900] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[901] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[902] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[903] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[904] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[905] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[906] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[907] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[908] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[909] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[910] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[911] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[912] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[913] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[914] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[915] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[916] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[917] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[918] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[919] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[920] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[921] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[922] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[923] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[924] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[925] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[926] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[927] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[928] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[929] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[930] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[931] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[932] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[933] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[934] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[935] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[936] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[937] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[938] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[939] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[940] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[941] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[942] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[943] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[944] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[945] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[946] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[947] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[948] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[949] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[950] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[951] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[952] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[953] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[954] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[955] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[956] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[957] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[958] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[959] = bs_data_in[0][3] & bs_data_in[1][2] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[960] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[961] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[962] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[963] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[964] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[965] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[966] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[967] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[968] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[969] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[970] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[971] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[972] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[973] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[974] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[975] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][0] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[976] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[977] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[978] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[979] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[980] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[981] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[982] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[983] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[984] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[985] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[986] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[987] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[988] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[989] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[990] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[991] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][1] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[992] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[993] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[994] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[995] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[996] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[997] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[998] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[999] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[1000] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[1001] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[1002] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[1003] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[1004] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[1005] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[1006] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[1007] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][2] & bs_data_in[3][3] & bs_data_in[4][3];
      assign bs_data_out[1008] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][0];
      assign bs_data_out[1009] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][1];
      assign bs_data_out[1010] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][2];
      assign bs_data_out[1011] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][0] & bs_data_in[4][3];
      assign bs_data_out[1012] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][0];
      assign bs_data_out[1013] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][1];
      assign bs_data_out[1014] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][2];
      assign bs_data_out[1015] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][1] & bs_data_in[4][3];
      assign bs_data_out[1016] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][0];
      assign bs_data_out[1017] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][1];
      assign bs_data_out[1018] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][2];
      assign bs_data_out[1019] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][2] & bs_data_in[4][3];
      assign bs_data_out[1020] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][0];
      assign bs_data_out[1021] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][1];
      assign bs_data_out[1022] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][2];
      assign bs_data_out[1023] = bs_data_in[0][3] & bs_data_in[1][3] & bs_data_in[2][3] & bs_data_in[3][3] & bs_data_in[4][3];

      par_acc_1024lanes  #(.WIDTH(WXIP1)) stoch2bin (
        .clk(clk),
        .rst(rst),                                               
        .data_in(bs_data_out),
        .countval(bin_data_out),
        .overflow(dummy_ov));

   end // if (NUM_INPUTS==5)
   
                                                            
    //FIXME 
	//assign done = sng_ov[NUM_INPUTS-1];
    assign done = sng_ov[NUM_INPUTS-1] | ~(|bs_data_in[NUM_INPUTS-1]);
    //assign done = sng_ov[NUM_INPUTS-1];
   
   


endmodule //ms_es_ordered_bs_by4_mul

