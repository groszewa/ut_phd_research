parameter DATA_WIDTH = 4;
parameter NUM_INPUTS = 2;
parameter WXIP1 = 9;
parameter MIN_CYC_DSC = 256;

